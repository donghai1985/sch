`ifndef PROJ_DEFINE_H
`define PROJ_DEFINE_H

//`define DEBUG_ILA
`define RDMA_MAX_SPEED
`define DDR4
`define RDMA_CHANNEL_1
`define RDMA_CHANNEL_2

`endif