// =================================================================================================
// Copyright(C) 2021 All rights reserved.
// =================================================================================================
//
// =================================================================================================
// File Name      : cmip_app_cnt.v
// Module         : cmip_app_cnt
// Function       : FPGA RTL Top module
// Type           : RTL
// -------------------------------------------------------------------------------------------------
// Update History :
// -------------------------------------------------------------------------------------------------
// Rev.Level  Date         Coded by         Contents
// 0.1.0      2020/02/03   NTEW)wang.qiuhua Create new
//
// =================================================================================================
// End Revision
// =================================================================================================

module cmip_app_cnt #(
    parameter WDTH = 16
)(
    input                          i_clk             ,//(i) 
    input                          i_rst_n           ,//(i) 
    input                          i_clr             ,//(i) 
    input                          i_vld             ,//(i) 
    output reg [WDTH-1:0]          o_cnt              //(o) 
);

// =================================================================================================
// RTL Body
// =================================================================================================
    reg     clr_d1;
    reg     clr_d2;


    always@(posedge i_clk)begin
        clr_d1 <= i_clr ;
        clr_d2 <= clr_d1;
    end



    always@(posedge i_clk or negedge i_rst_n)begin
       if(!i_rst_n)
          o_cnt <= {WDTH{1'b0}};
       else if(clr_d2)
          o_cnt <= {WDTH{1'b0}};
       else    if(i_vld)  
          o_cnt <= o_cnt +1'b1;
       else
          o_cnt <= o_cnt;
    end
          
          
          
    

endmodule





