`ifndef TDI_DEFINE_H
`define TDI_DEFINE_H

localparam TDI_0_width=35;		//35*64=2240
localparam TDI_0_width=37;		//37*64=2368

`endif