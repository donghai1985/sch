// =================================================================================================
// Copyright 2020 - 2030 (c) Inc. All rights reserved.
// =================================================================================================
//
// =================================================================================================
// File Name      : axidma_native.v
// Module         : axidma_native
// Type           : RTL
// -------------------------------------------------------------------------------------------------
// Update History :
// -------------------------------------------------------------------------------------------------
// Rev.Level  Date         Coded by         Contents
// 0.1.0      2022/12/14   NTEW)wang.qh     Create new
//
// =================================================================================================
// End Revision
// =================================================================================================

module axidma_inf #(
    parameter                               FIFO_DPTH       =  128         ,
    parameter                               DATA_WDTH       =  32          ,
    parameter                               ADDR_WDTH       =  32          ,
    parameter                               LEN_WDTH        =  32          
)(
    input                                   sys_clk                        ,//(i)
    input                                   sys_rst_n                      ,//(i)
    input                                   axi_clk                        ,//(i)
    input                                   axi_rst_n                      ,//(i)

    input                                   cfg_wsoft_rst                  ,//(i)
    input                                   cfg_wstart                     ,//(i)
    output                                  cfg_widle                      ,//(o)
    output            [LEN_WDTH -1:0]       cfg_wr_times                   ,//(o)
    input             [ADDR_WDTH-1:0]       cfg_base_waddr                 ,//(i)
    input             [LEN_WDTH -1:0]       cfg_wlen                       ,//(i)
    input             [7:0]                 cfg_wburst_len                 ,//(i)
    input                                   cfg_wirq_en                    ,//(i)
    input                                   cfg_wirq_clr                   ,//(i)
    output                                  wirq                           ,//(o)

    input                                   cfg_rsoft_rst                  ,//(i)
    input                                   cfg_rstart                     ,//(i)
    output                                  cfg_ridle                      ,//(i)
    output            [LEN_WDTH -1:0]       cfg_rd_times                   ,//(i)
    input             [ADDR_WDTH-1:0]       cfg_base_raddr                 ,//(i)
    input             [LEN_WDTH -1:0]       cfg_rlen                       ,//(i)
    input             [7:0]                 cfg_rburst_len                 ,//(i)
    input                                   cfg_rirq_en                    ,//(i)
    input                                   cfg_rirq_clr                   ,//(i)
    output                                  rirq                           ,//(o)

    // fifo wr ----> axi wr
    input                                   fifo_wr                        ,//(i)
    input             [DATA_WDTH-1:0]       fifo_din                       ,//(i)
    output                                  fifo_full                      ,//(o)
    // fifo rd <---- axi rd
    input                                   fifo_rd                        ,//(i)
    output            [DATA_WDTH-1:0]       fifo_dout                      ,//(i)
    output                                  fifo_empty                     ,//(o)

    output            [ADDR_WDTH-1:0]       m_axi_awaddr                   ,//(o)
    output            [ 1:0]                m_axi_awburst                  ,//(o)
    output            [ 3:0]                m_axi_awcache                  ,//(o)
    output            [ 3:0]                m_axi_awid                     ,//(o)
    output            [ 7:0]                m_axi_awlen                    ,//(o)
    output                                  m_axi_awlock                   ,//(o)
    output            [ 2:0]                m_axi_awprot                   ,//(o)
    output            [ 3:0]                m_axi_awqos                    ,//(o)
    output                                  m_axi_awvalid                  ,//(o)
    input                                   m_axi_awready                  ,//(i)
    output            [ 2:0]                m_axi_awsize                   ,//(o)
    output                                  m_axi_awuser                   ,//(o)
    input                                   m_axi_bvalid                   ,//(i)
    output                                  m_axi_bready                   ,//(o)
    input             [ 1:0]                m_axi_bresp                    ,//(i)
    input             [ 3:0]                m_axi_bid                      ,//(i)
    output                                  m_axi_wvalid                   ,//(o)
    input                                   m_axi_wready                   ,//(i)
    output            [DATA_WDTH/8-1:0]     m_axi_wstrb                    ,//(o)
    output            [DATA_WDTH-1:0]       m_axi_wdata                    ,//(o)
    output                                  m_axi_wlast                    ,//(o)

    output            [ADDR_WDTH-1:0]       m_axi_araddr                   ,//(o)
    output            [ 1:0]                m_axi_arburst                  ,//(o)
    output            [ 3:0]                m_axi_arcache                  ,//(o)
    output            [ 3:0]                m_axi_arid                     ,//(o)
    output            [ 7:0]                m_axi_arlen                    ,//(o)
    output                                  m_axi_arlock                   ,//(o)
    output            [ 2:0]                m_axi_arprot                   ,//(o)
    output            [ 3:0]                m_axi_arqos                    ,//(o)
    output                                  m_axi_arvalid                  ,//(o)
    input                                   m_axi_arready                  ,//(i)
    output            [ 2:0]                m_axi_arsize                   ,//(o)
    output                                  m_axi_aruser                   ,//(o)
    input             [DATA_WDTH-1:0]       m_axi_rdata                    ,//(i)
    input                                   m_axi_rvalid                   ,//(i)
    output                                  m_axi_rready                   ,//(o)
    input                                   m_axi_rlast                    ,//(i)
    input             [ 1:0]                m_axi_rresp                    ,//(i)
    input             [ 3:0]                m_axi_rid                       //(i)



);

    // -------------------------------------------------------------------------
    // Internal Parameter Definition
    // -------------------------------------------------------------------------    

    //---------------------------------------------------------------------
    // Defination of Internal Signals
    //---------------------------------------------------------------------
    // wire                                cfg_wsoft_rst                      ;
    // wire                                cfg_wstart                         ;
    // wire                                cfg_widle                          ;
    // wire          [LEN_WDTH -1:0]       cfg_wr_times                       ;
    // wire          [ADDR_WDTH-1:0]       cfg_base_waddr                     ;
    // wire          [LEN_WDTH -1:0]       cfg_wlen                           ;
    // wire          [7:0]                 cfg_wburst_len                     ;
    // wire                                cfg_wirq_en                        ;
    // wire                                cfg_wirq_clr                       ;

    wire                                wstart_vld                         ;
    wire                                wstart_rdy                         ;
    wire          [ADDR_WDTH-1:0]       waddr                              ;
    wire          [7:0]                 wburst_len                         ;

    // wire                                cfg_rsoft_rst                      ;
    // wire                                cfg_rstart                         ;
    // wire                                cfg_ridle                          ;
    // wire          [LEN_WDTH -1:0]       cfg_rd_times                       ;
    // wire          [ADDR_WDTH-1:0]       cfg_base_raddr                     ;
    // wire          [LEN_WDTH -1:0]       cfg_rlen                           ;
    // wire          [7:0]                 cfg_rburst_len                     ;
    // wire                                cfg_rirq_en                        ;
    // wire                                cfg_rirq_clr                       ;

    wire                                rstart_vld                         ;
    wire                                rstart_rdy                         ;
    wire          [ADDR_WDTH-1:0]       raddr                              ;
    wire          [7:0]                 rburst_len                         ;


    // -------------------------------------------------------------------------
    // output
    // -------------------------------------------------------------------------


// =================================================================================================
// RTL Body
// =================================================================================================
    axidma_wr_fsm #(
        .LEN_WDTH                       (LEN_WDTH                ),
        .DATA_WDTH                      (DATA_WDTH               ),
        .ADDR_WDTH                      (ADDR_WDTH               )
    )u_axidma_wr_fsm(                   
        .sys_clk                        (axi_clk                 ),//(i)
        .sys_rst_n                      (axi_rst_n               ),//(i)
        .cfg_wburst_len                 (cfg_wburst_len          ),//(i)
        .cfg_wsoft_rst                  (cfg_wsoft_rst           ),//(i)
        .cfg_wstart                     (cfg_wstart              ),//(i)
        .cfg_waddr                      (cfg_base_waddr          ),//(i)
        .cfg_wlen                       (cfg_wlen                ),//(i)
        .cfg_widle                      (cfg_widle               ),//(o)
        .cfg_wr_times                   (cfg_wr_times            ),//(o)
        .cfg_wirq_en                    (cfg_wirq_en             ),//(i)
        .cfg_wirq_clr                   (cfg_wirq_clr            ),//(i)
        .wirq                           (wirq                    ),//(o)

        .wstart_vld                     (wstart_vld              ),//(i)
        .wstart_rdy                     (wstart_rdy              ),//(o)
        .waddr                          (waddr                   ),//(i)
        .wburst_len                     (wburst_len              ) //(i)
    );


    axidma_rd_fsm #(
        .LEN_WDTH                       (LEN_WDTH                ),
        .DATA_WDTH                      (DATA_WDTH               ),
        .ADDR_WDTH                      (ADDR_WDTH               )
    )u_axidma_rd_fsm(                                                   
        .sys_clk                        (axi_clk                 ),//(i)
        .sys_rst_n                      (axi_rst_n               ),//(i)
        .cfg_rburst_len                 (cfg_rburst_len          ),//(i)
        .cfg_rsoft_rst                  (cfg_rsoft_rst           ),//(i)
        .cfg_rstart                     (cfg_rstart              ),//(i)
        .cfg_raddr                      (cfg_base_raddr          ),//(i)
        .cfg_rlen                       (cfg_rlen                ),//(i)
        .cfg_ridle                      (cfg_ridle               ),//(o)
        .cfg_rd_times                   (cfg_rd_times            ),//(o)
        .cfg_rirq_en                    (cfg_rirq_en             ),//(i)
        .cfg_rirq_clr                   (cfg_rirq_clr            ),//(i)
        .rirq                           (rirq                    ),//(o)

        .rstart_vld                     (rstart_vld              ),//(i)
        .rstart_rdy                     (rstart_rdy              ),//(o)
        .raddr                          (raddr                   ),//(i)
        .rburst_len                     (rburst_len              ) //(i)
    );


    fifo2axi_native #(
        .FIFO_DPTH                      (FIFO_DPTH        ),
        .DATA_WDTH                      (DATA_WDTH        ),
        .ADDR_WDTH                      (ADDR_WDTH        )
    )u_fifo2axi_native(                                          
        .sys_clk                        (sys_clk          ),//(i)
        .sys_rst_n                      (sys_rst_n        ),//(i)
        .axi_clk                        (axi_clk          ),//(i)
        .axi_rst_n                      (axi_rst_n        ),//(i)
        .fifo_wr                        (fifo_wr          ),//(i)
        .fifo_din                       (fifo_din         ),//(i)
        .fifo_full                      (fifo_full        ),//(o)
        .wsoft_rst                      (cfg_wsoft_rst    ),//(i)
        .wstart_vld                     (wstart_vld       ),//(i)
        .wstart_rdy                     (wstart_rdy       ),//(o)
        .waddr                          (waddr            ),//(i)
        .wburst_len                     (wburst_len       ),//(i)

        .m_axi_awaddr                   (m_axi_awaddr     ),//(o)
        .m_axi_awburst                  (m_axi_awburst    ),//(o)
        .m_axi_awcache                  (m_axi_awcache    ),//(o)
        .m_axi_awid                     (m_axi_awid       ),//(o)
        .m_axi_awlen                    (m_axi_awlen      ),//(o)
        .m_axi_awlock                   (m_axi_awlock     ),//(o)
        .m_axi_awprot                   (m_axi_awprot     ),//(o)
        .m_axi_awqos                    (m_axi_awqos      ),//(o)
        .m_axi_awvalid                  (m_axi_awvalid    ),//(o)
        .m_axi_awready                  (m_axi_awready    ),//(i)
        .m_axi_awsize                   (m_axi_awsize     ),//(o)
        .m_axi_awuser                   (m_axi_awuser     ),//(o)
        .m_axi_bvalid                   (m_axi_bvalid     ),//(i)
        .m_axi_bready                   (m_axi_bready     ),//(o)
        .m_axi_bresp                    (m_axi_bresp      ),//(i)
        .m_axi_bid                      (m_axi_bid        ),//(i)
        .m_axi_wvalid                   (m_axi_wvalid     ),//(o)
        .m_axi_wready                   (m_axi_wready     ),//(i)
        .m_axi_wstrb                    (m_axi_wstrb      ),//(o)
        .m_axi_wdata                    (m_axi_wdata      ),//(o)
        .m_axi_wlast                    (m_axi_wlast      ),//(o)

        .fifo_rd                        (fifo_rd          ),//(i)
        .fifo_dout                      (fifo_dout        ),//(i)
        .fifo_empty                     (fifo_empty       ),//(o)
        .rsoft_rst                      (cfg_rsoft_rst    ),//(i)
        .rstart_vld                     (rstart_vld       ),//(i)
        .rstart_rdy                     (rstart_rdy       ),//(o)
        .raddr                          (raddr            ),//(i)
        .rburst_len                     (rburst_len       ),//(i)

        .m_axi_araddr                   (m_axi_araddr     ),//(o)
        .m_axi_arburst                  (m_axi_arburst    ),//(o)
        .m_axi_arcache                  (m_axi_arcache    ),//(o)
        .m_axi_arid                     (m_axi_arid       ),//(o)
        .m_axi_arlen                    (m_axi_arlen      ),//(o)
        .m_axi_arlock                   (m_axi_arlock     ),//(o)
        .m_axi_arprot                   (m_axi_arprot     ),//(o)
        .m_axi_arqos                    (m_axi_arqos      ),//(o)
        .m_axi_arvalid                  (m_axi_arvalid    ),//(o)
        .m_axi_arready                  (m_axi_arready    ),//(i)
        .m_axi_arsize                   (m_axi_arsize     ),//(o)
        .m_axi_aruser                   (m_axi_aruser     ),//(o)
        .m_axi_rdata                    (m_axi_rdata      ),//(i)
        .m_axi_rvalid                   (m_axi_rvalid     ),//(i)
        .m_axi_rready                   (m_axi_rready     ),//(o)
        .m_axi_rlast                    (m_axi_rlast      ),//(i)
        .m_axi_rresp                    (m_axi_rresp      ),//(i)
        .m_axi_rid                      (m_axi_rid        ) //(i)
    );































endmodule





